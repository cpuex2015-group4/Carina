--bclt
--bclf
--lw.s
--sw.s

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

library work;
use work.p_type.all;


entity arith_core is
  clk:in std_logic;
  IO_recv_data
end arith_core;
